`include  "add_overflow_class.sv"
`timescale 1ps / 1ps
module test;
reg  clk;
reg  rst_n;
reg  enable;
reg  [1:0]rounding;
reg  [2:0]operation;
reg  [63:0]operand_a;
reg  [63:0]operand_b;
wire  [63:0]out;
wire  ready;
wire  underflow;
wire  overflow;
wire  inexact;
wire  exception;
wire  invalid;
fpu ins1 (
.clk(clk),
.rst_n(rst_n),
.enable(enable),
.rounding(rounding),
.operation(operation),
.operand_a(operand_a),
.operand_b(operand_b),
.out(out),
.ready(ready),
.underflow(underflow),
.overflow(overflow),
.inexact(inexact),
.exception(exception),
.invalid(invalid)
);
packet0  p0;
packet1  p1;
packet2  p2;
packet3  p3;
packet4  p4;
packet5  p5;
packet6  p6;
packet7  p7;
packet8  p8;
packet9  p9;
packet10  p10;
packet11  p11;
packet12  p12;
packet13  p13;
packet14  p14;
packet15  p15;
initial
begin
p0=new();
p1=new();
p2=new();
p3=new();
p4=new();
p5=new();
p6=new();
p7=new();
p8=new();
p9=new();
p10=new();
p11=new();
p12=new();
p13=new();
p14=new();
p15=new();
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p0.constraint_mode(0);
p0.c0.constraint_mode(1);
assert(p0.randomize());
rst_n=p0.rst_n;
enable=p0.enable;
rounding=p0.rounding;
operation=p0.operation;
operand_a=p0.operand_a;
operand_b=p0.operand_b;
p0.out=out;
p0.ready=ready;
p0.underflow=underflow;
p0.overflow=overflow;
p0.inexact=inexact;
p0.exception=exception;
p0.invalid=invalid;
#20000;
p0.constraint_mode(0);
p0.c1.constraint_mode(1);
assert(p0.randomize(enable));
rst_n=p0.rst_n;
enable=p0.enable;
rounding=p0.rounding;
operation=p0.operation;
operand_a=p0.operand_a;
operand_b=p0.operand_b;
p0.out=out;
p0.ready=ready;
p0.underflow=underflow;
p0.overflow=overflow;
p0.inexact=inexact;
p0.exception=exception;
p0.invalid=invalid;
#800000;
p0.constraint_mode(0);
p0.c2.constraint_mode(1);
assert(p0.randomize(overflow,enable,operand_a,operand_b));
rst_n=p0.rst_n;
enable=p0.enable;
rounding=p0.rounding;
operation=p0.operation;
operand_a=p0.operand_a;
operand_b=p0.operand_b;
p0.out=out;
p0.ready=ready;
p0.underflow=underflow;
p0.overflow=overflow;
p0.inexact=inexact;
p0.exception=exception;
p0.invalid=invalid;
#20000;
p0.constraint_mode(0);
p0.c3.constraint_mode(1);
assert(p0.randomize(enable));
rst_n=p0.rst_n;
enable=p0.enable;
rounding=p0.rounding;
operation=p0.operation;
operand_a=p0.operand_a;
operand_b=p0.operand_b;
p0.out=out;
p0.ready=ready;
p0.underflow=underflow;
p0.overflow=overflow;
p0.inexact=inexact;
p0.exception=exception;
p0.invalid=invalid;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p1.constraint_mode(0);
p1.c0.constraint_mode(1);
assert(p1.randomize());
rst_n=p1.rst_n;
enable=p1.enable;
rounding=p1.rounding;
operation=p1.operation;
operand_a=p1.operand_a;
operand_b=p1.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p1.constraint_mode(0);
p1.c1.constraint_mode(1);
assert(p1.randomize(enable));
rst_n=p1.rst_n;
enable=p1.enable;
rounding=p1.rounding;
operation=p1.operation;
operand_a=p1.operand_a;
operand_b=p1.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p1.constraint_mode(0);
p1.c2.constraint_mode(1);
assert(p1.randomize(overflow,enable,operand_a,operand_b));
rst_n=p1.rst_n;
enable=p1.enable;
rounding=p1.rounding;
operation=p1.operation;
operand_a=p1.operand_a;
operand_b=p1.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p1.constraint_mode(0);
p1.c3.constraint_mode(1);
assert(p1.randomize(enable));
rst_n=p1.rst_n;
enable=p1.enable;
rounding=p1.rounding;
operation=p1.operation;
operand_a=p1.operand_a;
operand_b=p1.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p2.constraint_mode(0);
p2.c0.constraint_mode(1);
assert(p2.randomize());
rst_n=p2.rst_n;
enable=p2.enable;
rounding=p2.rounding;
operation=p2.operation;
operand_a=p2.operand_a;
operand_b=p2.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p2.constraint_mode(0);
p2.c1.constraint_mode(1);
assert(p2.randomize(enable));
rst_n=p2.rst_n;
enable=p2.enable;
rounding=p2.rounding;
operation=p2.operation;
operand_a=p2.operand_a;
operand_b=p2.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p2.constraint_mode(0);
p2.c2.constraint_mode(1);
assert(p2.randomize(overflow,enable,operand_a,operand_b));
rst_n=p2.rst_n;
enable=p2.enable;
rounding=p2.rounding;
operation=p2.operation;
operand_a=p2.operand_a;
operand_b=p2.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p2.constraint_mode(0);
p2.c3.constraint_mode(1);
assert(p2.randomize(enable));
rst_n=p2.rst_n;
enable=p2.enable;
rounding=p2.rounding;
operation=p2.operation;
operand_a=p2.operand_a;
operand_b=p2.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p3.constraint_mode(0);
p3.c0.constraint_mode(1);
assert(p3.randomize());
rst_n=p3.rst_n;
enable=p3.enable;
rounding=p3.rounding;
operation=p3.operation;
operand_a=p3.operand_a;
operand_b=p3.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p3.constraint_mode(0);
p3.c1.constraint_mode(1);
assert(p3.randomize(enable));
rst_n=p3.rst_n;
enable=p3.enable;
rounding=p3.rounding;
operation=p3.operation;
operand_a=p3.operand_a;
operand_b=p3.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p3.constraint_mode(0);
p3.c2.constraint_mode(1);
assert(p3.randomize(overflow,enable,operand_a,operand_b));
rst_n=p3.rst_n;
enable=p3.enable;
rounding=p3.rounding;
operation=p3.operation;
operand_a=p3.operand_a;
operand_b=p3.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p3.constraint_mode(0);
p3.c3.constraint_mode(1);
assert(p3.randomize(enable));
rst_n=p3.rst_n;
enable=p3.enable;
rounding=p3.rounding;
operation=p3.operation;
operand_a=p3.operand_a;
operand_b=p3.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p4.constraint_mode(0);
p4.c0.constraint_mode(1);
assert(p4.randomize());
rst_n=p4.rst_n;
enable=p4.enable;
rounding=p4.rounding;
operation=p4.operation;
operand_a=p4.operand_a;
operand_b=p4.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p4.constraint_mode(0);
p4.c1.constraint_mode(1);
assert(p4.randomize(enable));
rst_n=p4.rst_n;
enable=p4.enable;
rounding=p4.rounding;
operation=p4.operation;
operand_a=p4.operand_a;
operand_b=p4.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p4.constraint_mode(0);
p4.c2.constraint_mode(1);
assert(p4.randomize(overflow,enable,operand_a,operand_b));
rst_n=p4.rst_n;
enable=p4.enable;
rounding=p4.rounding;
operation=p4.operation;
operand_a=p4.operand_a;
operand_b=p4.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p4.constraint_mode(0);
p4.c3.constraint_mode(1);
assert(p4.randomize(enable));
rst_n=p4.rst_n;
enable=p4.enable;
rounding=p4.rounding;
operation=p4.operation;
operand_a=p4.operand_a;
operand_b=p4.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p5.constraint_mode(0);
p5.c0.constraint_mode(1);
assert(p5.randomize());
rst_n=p5.rst_n;
enable=p5.enable;
rounding=p5.rounding;
operation=p5.operation;
operand_a=p5.operand_a;
operand_b=p5.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p5.constraint_mode(0);
p5.c1.constraint_mode(1);
assert(p5.randomize(enable));
rst_n=p5.rst_n;
enable=p5.enable;
rounding=p5.rounding;
operation=p5.operation;
operand_a=p5.operand_a;
operand_b=p5.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p5.constraint_mode(0);
p5.c2.constraint_mode(1);
assert(p5.randomize(overflow,enable,operand_a,operand_b));
rst_n=p5.rst_n;
enable=p5.enable;
rounding=p5.rounding;
operation=p5.operation;
operand_a=p5.operand_a;
operand_b=p5.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p5.constraint_mode(0);
p5.c3.constraint_mode(1);
assert(p5.randomize(enable));
rst_n=p5.rst_n;
enable=p5.enable;
rounding=p5.rounding;
operation=p5.operation;
operand_a=p5.operand_a;
operand_b=p5.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p6.constraint_mode(0);
p6.c0.constraint_mode(1);
assert(p6.randomize());
rst_n=p6.rst_n;
enable=p6.enable;
rounding=p6.rounding;
operation=p6.operation;
operand_a=p6.operand_a;
operand_b=p6.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p6.constraint_mode(0);
p6.c1.constraint_mode(1);
assert(p6.randomize(enable));
rst_n=p6.rst_n;
enable=p6.enable;
rounding=p6.rounding;
operation=p6.operation;
operand_a=p6.operand_a;
operand_b=p6.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p6.constraint_mode(0);
p6.c2.constraint_mode(1);
assert(p6.randomize(overflow,enable,operand_a,operand_b));
rst_n=p6.rst_n;
enable=p6.enable;
rounding=p6.rounding;
operation=p6.operation;
operand_a=p6.operand_a;
operand_b=p6.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p6.constraint_mode(0);
p6.c3.constraint_mode(1);
assert(p6.randomize(enable));
rst_n=p6.rst_n;
enable=p6.enable;
rounding=p6.rounding;
operation=p6.operation;
operand_a=p6.operand_a;
operand_b=p6.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p7.constraint_mode(0);
p7.c0.constraint_mode(1);
assert(p7.randomize());
rst_n=p7.rst_n;
enable=p7.enable;
rounding=p7.rounding;
operation=p7.operation;
operand_a=p7.operand_a;
operand_b=p7.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p7.constraint_mode(0);
p7.c1.constraint_mode(1);
assert(p7.randomize(enable));
rst_n=p7.rst_n;
enable=p7.enable;
rounding=p7.rounding;
operation=p7.operation;
operand_a=p7.operand_a;
operand_b=p7.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p7.constraint_mode(0);
p7.c2.constraint_mode(1);
assert(p7.randomize(overflow,enable,operand_a,operand_b));
rst_n=p7.rst_n;
enable=p7.enable;
rounding=p7.rounding;
operation=p7.operation;
operand_a=p7.operand_a;
operand_b=p7.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p7.constraint_mode(0);
p7.c3.constraint_mode(1);
assert(p7.randomize(enable));
rst_n=p7.rst_n;
enable=p7.enable;
rounding=p7.rounding;
operation=p7.operation;
operand_a=p7.operand_a;
operand_b=p7.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p8.constraint_mode(0);
p8.c0.constraint_mode(1);
assert(p8.randomize());
rst_n=p8.rst_n;
enable=p8.enable;
rounding=p8.rounding;
operation=p8.operation;
operand_a=p8.operand_a;
operand_b=p8.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p8.constraint_mode(0);
p8.c1.constraint_mode(1);
assert(p8.randomize(enable));
rst_n=p8.rst_n;
enable=p8.enable;
rounding=p8.rounding;
operation=p8.operation;
operand_a=p8.operand_a;
operand_b=p8.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p8.constraint_mode(0);
p8.c2.constraint_mode(1);
assert(p8.randomize(overflow,enable,operand_a,operand_b));
rst_n=p8.rst_n;
enable=p8.enable;
rounding=p8.rounding;
operation=p8.operation;
operand_a=p8.operand_a;
operand_b=p8.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p8.constraint_mode(0);
p8.c3.constraint_mode(1);
assert(p8.randomize(enable));
rst_n=p8.rst_n;
enable=p8.enable;
rounding=p8.rounding;
operation=p8.operation;
operand_a=p8.operand_a;
operand_b=p8.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p9.constraint_mode(0);
p9.c0.constraint_mode(1);
assert(p9.randomize());
rst_n=p9.rst_n;
enable=p9.enable;
rounding=p9.rounding;
operation=p9.operation;
operand_a=p9.operand_a;
operand_b=p9.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p9.constraint_mode(0);
p9.c1.constraint_mode(1);
assert(p9.randomize(enable));
rst_n=p9.rst_n;
enable=p9.enable;
rounding=p9.rounding;
operation=p9.operation;
operand_a=p9.operand_a;
operand_b=p9.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p9.constraint_mode(0);
p9.c2.constraint_mode(1);
assert(p9.randomize(overflow,enable,operand_a,operand_b));
rst_n=p9.rst_n;
enable=p9.enable;
rounding=p9.rounding;
operation=p9.operation;
operand_a=p9.operand_a;
operand_b=p9.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p9.constraint_mode(0);
p9.c3.constraint_mode(1);
assert(p9.randomize(enable));
rst_n=p9.rst_n;
enable=p9.enable;
rounding=p9.rounding;
operation=p9.operation;
operand_a=p9.operand_a;
operand_b=p9.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p10.constraint_mode(0);
p10.c0.constraint_mode(1);
assert(p10.randomize());
rst_n=p10.rst_n;
enable=p10.enable;
rounding=p10.rounding;
operation=p10.operation;
operand_a=p10.operand_a;
operand_b=p10.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p10.constraint_mode(0);
p10.c1.constraint_mode(1);
assert(p10.randomize(enable));
rst_n=p10.rst_n;
enable=p10.enable;
rounding=p10.rounding;
operation=p10.operation;
operand_a=p10.operand_a;
operand_b=p10.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p10.constraint_mode(0);
p10.c2.constraint_mode(1);
assert(p10.randomize(overflow,enable,operand_a,operand_b));
rst_n=p10.rst_n;
enable=p10.enable;
rounding=p10.rounding;
operation=p10.operation;
operand_a=p10.operand_a;
operand_b=p10.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p10.constraint_mode(0);
p10.c3.constraint_mode(1);
assert(p10.randomize(enable));
rst_n=p10.rst_n;
enable=p10.enable;
rounding=p10.rounding;
operation=p10.operation;
operand_a=p10.operand_a;
operand_b=p10.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p11.constraint_mode(0);
p11.c0.constraint_mode(1);
assert(p11.randomize());
rst_n=p11.rst_n;
enable=p11.enable;
rounding=p11.rounding;
operation=p11.operation;
operand_a=p11.operand_a;
operand_b=p11.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p11.constraint_mode(0);
p11.c1.constraint_mode(1);
assert(p11.randomize(enable));
rst_n=p11.rst_n;
enable=p11.enable;
rounding=p11.rounding;
operation=p11.operation;
operand_a=p11.operand_a;
operand_b=p11.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p11.constraint_mode(0);
p11.c2.constraint_mode(1);
assert(p11.randomize(overflow,enable,operand_a,operand_b));
rst_n=p11.rst_n;
enable=p11.enable;
rounding=p11.rounding;
operation=p11.operation;
operand_a=p11.operand_a;
operand_b=p11.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p11.constraint_mode(0);
p11.c3.constraint_mode(1);
assert(p11.randomize(enable));
rst_n=p11.rst_n;
enable=p11.enable;
rounding=p11.rounding;
operation=p11.operation;
operand_a=p11.operand_a;
operand_b=p11.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p12.constraint_mode(0);
p12.c0.constraint_mode(1);
assert(p12.randomize());
rst_n=p12.rst_n;
enable=p12.enable;
rounding=p12.rounding;
operation=p12.operation;
operand_a=p12.operand_a;
operand_b=p12.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p12.constraint_mode(0);
p12.c1.constraint_mode(1);
assert(p12.randomize(enable));
rst_n=p12.rst_n;
enable=p12.enable;
rounding=p12.rounding;
operation=p12.operation;
operand_a=p12.operand_a;
operand_b=p12.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p12.constraint_mode(0);
p12.c2.constraint_mode(1);
assert(p12.randomize(overflow,enable,operand_a,operand_b));
rst_n=p12.rst_n;
enable=p12.enable;
rounding=p12.rounding;
operation=p12.operation;
operand_a=p12.operand_a;
operand_b=p12.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p12.constraint_mode(0);
p12.c3.constraint_mode(1);
assert(p12.randomize(enable));
rst_n=p12.rst_n;
enable=p12.enable;
rounding=p12.rounding;
operation=p12.operation;
operand_a=p12.operand_a;
operand_b=p12.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p13.constraint_mode(0);
p13.c0.constraint_mode(1);
assert(p13.randomize());
rst_n=p13.rst_n;
enable=p13.enable;
rounding=p13.rounding;
operation=p13.operation;
operand_a=p13.operand_a;
operand_b=p13.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p13.constraint_mode(0);
p13.c1.constraint_mode(1);
assert(p13.randomize(enable));
rst_n=p13.rst_n;
enable=p13.enable;
rounding=p13.rounding;
operation=p13.operation;
operand_a=p13.operand_a;
operand_b=p13.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p13.constraint_mode(0);
p13.c2.constraint_mode(1);
assert(p13.randomize(overflow,enable,operand_a,operand_b));
rst_n=p13.rst_n;
enable=p13.enable;
rounding=p13.rounding;
operation=p13.operation;
operand_a=p13.operand_a;
operand_b=p13.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p13.constraint_mode(0);
p13.c3.constraint_mode(1);
assert(p13.randomize(enable));
rst_n=p13.rst_n;
enable=p13.enable;
rounding=p13.rounding;
operation=p13.operation;
operand_a=p13.operand_a;
operand_b=p13.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p14.constraint_mode(0);
p14.c0.constraint_mode(1);
assert(p14.randomize());
rst_n=p14.rst_n;
enable=p14.enable;
rounding=p14.rounding;
operation=p14.operation;
operand_a=p14.operand_a;
operand_b=p14.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p14.constraint_mode(0);
p14.c1.constraint_mode(1);
assert(p14.randomize(enable));
rst_n=p14.rst_n;
enable=p14.enable;
rounding=p14.rounding;
operation=p14.operation;
operand_a=p14.operand_a;
operand_b=p14.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p14.constraint_mode(0);
p14.c2.constraint_mode(1);
assert(p14.randomize(overflow,enable,operand_a,operand_b));
rst_n=p14.rst_n;
enable=p14.enable;
rounding=p14.rounding;
operation=p14.operation;
operand_a=p14.operand_a;
operand_b=p14.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p14.constraint_mode(0);
p14.c3.constraint_mode(1);
assert(p14.randomize(enable));
rst_n=p14.rst_n;
enable=p14.enable;
rounding=p14.rounding;
operation=p14.operation;
operand_a=p14.operand_a;
operand_b=p14.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
#0
rst_n = 1'b1;
# 20000;
repeat(100)
begin

p15.constraint_mode(0);
p15.c0.constraint_mode(1);
assert(p15.randomize());
rst_n=p15.rst_n;
enable=p15.enable;
rounding=p15.rounding;
operation=p15.operation;
operand_a=p15.operand_a;
operand_b=p15.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p15.constraint_mode(0);
p15.c1.constraint_mode(1);
assert(p15.randomize(enable));
rst_n=p15.rst_n;
enable=p15.enable;
rounding=p15.rounding;
operation=p15.operation;
operand_a=p15.operand_a;
operand_b=p15.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#800000;
p15.constraint_mode(0);
p15.c2.constraint_mode(1);
assert(p15.randomize(overflow,enable,operand_a,operand_b));
rst_n=p15.rst_n;
enable=p15.enable;
rounding=p15.rounding;
operation=p15.operation;
operand_a=p15.operand_a;
operand_b=p15.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
#20000;
p15.constraint_mode(0);
p15.c3.constraint_mode(1);
assert(p15.randomize(enable));
rst_n=p15.rst_n;
enable=p15.enable;
rounding=p15.rounding;
operation=p15.operation;
operand_a=p15.operand_a;
operand_b=p15.operand_b;
# 800000;
$display("rst_n=%b",rst_n);
$display("enable=%b",enable);
$display("rounding=%b",rounding);
$display("operation=%b",operation);
$display("operand_a=%b",operand_a);
$display("operand_b=%b",operand_b);
$display("out=%b",out);
$display("ready=%b",ready);
$display("underflow=%b",underflow);
$display("overflow=%b",overflow);
$display("inexact=%b",inexact);
$display("exception=%b",exception);
$display("invalid=%b",invalid);
end
$finish;
end
always
begin : CLOCK_clk
clk = 1'b0;
#5000;
clk = 1'b1;
#5000;
end
endmodule
